/*	 ___________________________________________
	|											|
	|			   _    ____  _   _ 			|
	|			  / \  |  _ \| | | |			|
	|			 / _ \ | |_) | | | |			|
	|			/ ___ \|  __/| |_| |			|
	|		   /_/   \_|_|    \___/ 			|
	|		The Audio Processing Unit			|
	|											|
	|___________________________________________|
	
	
	The NES APU has 5 programmable sound generators. The base frequency used to generate all sounds is the CPU frequency







*/
`define BYTE reg[7:0]

module apu();
	BYTE cRegs[0:21];		/*
								
							*/
	
endmodule